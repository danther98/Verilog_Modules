module CLA16_tb();
reg [15:0] X;
reg [15:0] Y;
reg Cin;
wire [15:0] S;
wire Co;
CLA16 CLA16_1(.S(S),.Co(Co),.X(X),.Y(Y),.Cin(Cin));
initial begin
X = 16'b0;
Y = 16'b0;
Cin = 0;
#100;
X=16'b0000000000000001;
Y=16'b0000000000000001;
Cin=0;
#50;
X=16'b0000000000000010;
Y=16'b0000000000000010;
Cin=0;
#50;
X=16'b0000000000000011;
Y=16'b0000000000000011;
Cin=0;
#50;
X=16'b0000000000000100;
Y=16'b0000000000000100;
Cin=0;
#50;
X=16'b0000000000000101;
Y=16'b0000000000000101;
Cin=0;
#50;
X=16'b0000000000000110;
Y=16'b0000000000000110;
Cin=0;
#50;
X=16'b0000000000000111;
Y=16'b0000000000000111;
Cin=0;
#50;
X=16'b0000000000001000;
Y=16'b0000000000001000;
Cin=0;
#50;
X=16'b0000000000001001;
Y=16'b0000000000001001;
Cin=0;
#50;
X=16'b0000000000001010;
Y=16'b0000000000001010;
Cin=0;
#50;
X=16'b0000000000001011;
Y=16'b0000000000001011;
Cin=0;
#50;
Cin=1;
#100;



end


endmodule


